module riscv_hart
(
	input	wire		clk,
	input	wire		rst,

	output	wire		imem_addr_valid,
	output	wire	[31:0]	imem_addr,
	input	wire		imem_data_ready,
	input	wire	[31:0]	imem_data,

	output	wire	[2:0]	dmem_op,
	output	wire		dmem_addr_valid,
	output	wire	[31:0]	dmem_addr,
	input	wire		dmem_read_data_ready,
	input	wire	[31:0]	dmem_read_data,
	output	wire		dmem_write_data_valid,
	output	wire	[31:0]	dmem_write_data,

	input	wire		hardware_irq,
	input	wire		timer_irq
);

integer i;

wire		illegal_instruction;
wire		breakpoint;
wire		ecall;
wire		trap;
wire		mret;
wire		wfi;
wire	[31:0]	trap_target;
wire	[31:0]	mret_target;
wire	[31:0]	nextpc;
wire	[4:0]	rs1;
wire	[4:0]	rs2;
wire	[11:0]	csr;
wire	[4095:0]	csr_;
wire	[31:0]	csr_value;
wire		jump;
wire	[31:0]	jump_target;
wire	[4:0]	rd;
wire	[31:0]	csr_wb;
wire	[31:0]	irf_wb;

// Main operation registers

reg	[31:0]	pc;
reg	[31:0]	instr;
reg	[31:0]	irf	[0:31];


// Initialize regs

initial
begin
	pc = -4;
	instr = 32'h13;

	for (i = 0; i < 32; i++)
	begin
		irf[i] = 0;
	end
end

riscv_control control
(
	.clk(clk),
	.rst(rst),

	// CSR read/write port
	.csr(csr),
	.csr_(csr_),
	.csr_value(csr_value),
	.csr_wb(csr_wb),

	// Memory access monitoring port
	.pc(pc),
	.imem_data_ready(imem_data_ready),
	.dmem_op(dmem_op),
	.addr(dmem_addr),

	// Inline event port
	.illegal_instruction(illegal_instruction),
	.breakpoint(breakpoint),
	.ecall(ecall),
	.mret(mret),
	.wfi(wfi),

	// Interrupt port
	.hardware_irq(hardware_irq),
	.timer_irq(timer_irq),

	// Trap port
	.trap(trap),
	.trap_target(trap_target),
	.mret_target(mret_target)
);


// Fetch logic

assign nextpc =	rst ?				0 :
		trap ?				trap_target :
		wfi ?				pc :
		mret ?				mret_target :
		jump ?				jump_target :
						pc + 4;

assign imem_addr_valid = 1;
assign imem_addr = nextpc;

always @(posedge clk, posedge rst)
begin
	if (rst)
	begin
		pc <= -4;
		instr <= 32'h13;
	end else if (imem_data_ready & (dmem_addr_valid ? dmem_read_data_ready : 1))
	begin
		pc <= nextpc;
		instr <= imem_data;
	end
end


riscv_datapath datapath
(
	.clk(clk),

	// instruction/pc input
	.pc(pc),
	.instr(instr),

	// exception detection port
	.illegal_instruction(illegal_instruction),
	.breakpoint(breakpoint),
	.ecall(ecall),
	.mret(mret),
	.wfi(wfi),

	// irf read port
	.rs1(rs1),
	.rs2(rs2),
	.rs1_value(irf[rs1]),
	.rs2_value(irf[rs2]),

	// csr read/write port
	.csr(csr),
	.csr_(csr_),
	.csr_value(csr_value),
	.csr_wb(csr_wb),

	// jump port
	.jump(jump),
	.jump_target(jump_target),

	// memory access port 
	.is_mem_op(dmem_addr_valid),
	.is_store(dmem_write_data_valid),
	.mem_op(dmem_op),
	.mem_addr(dmem_addr),
	.mem_load_data(dmem_read_data),
	.mem_store_data(dmem_write_data),

	// irf writeback port 
	.rd(rd),
	.irf_wb(irf_wb)
);

// Writeback

always @(posedge clk, posedge rst)
begin
	if (rst)
	begin
		for (i = 0; i < 32; i++)
		begin
			irf[i] <= 32'b0;
		end
	end else if ((rd != 5'b0) & imem_data_ready)
	begin
		irf[rd] <= irf_wb;
	end
end

endmodule
